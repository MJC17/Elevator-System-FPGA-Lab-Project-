// Module to generate a slower clock signal (CLK_out) from a faster input clock (CLK_in)
module Adjust_Clk( CLK_in, CLK_out);
    input CLK_in;  // Input clock signal (50 MHz)
    output CLK_out; // Output slower clock signal
    reg [26:0] count = 0; // 27-bit counter used to divide the clock frequency

    // Always block triggered on every rising edge of the input clock (CLK_in)
    always @(posedge CLK_in) begin
        count <= count + 1'b1;  // Increment counter by 1 on each rising edge of CLK_in
    end

    // Assign the 23rd bit of the counter to the output clock (CLK_out), 
    // generating a slower clock (approximately 3 Hz)
    assign CLK_out = count[23]; // The slower clock derived from the 23rd bit of the counter
endmodule

// Main module representing the Elevator System
module LabElevatorProject(
    input CLK_50MHz, floorBtn1, floorBtn2, floorBtn3, // Floor buttons to select desired floor
    floorSwitch1, floorSwitch2, floorSwitch3, // Reed switches to detect the current elevator position
    output reg LEDA, LEDB, LEDC, LEDD, LEDE, LEDF, LEDG, LED0, LED1, LED2, UpPin, DownPin
);
    // Internal registers to hold the state of the elevator system
    reg [6:0] LevelLights = 7'b1111111;  // Default level, all LEDs off
    reg [1:0] SelectedLevel = 2'b00;  // Initialize the selected floor to floor 0 (2 bits)
    reg [1:0] CurrentLevel = 2'b00;   // Initialize the current floor to floor 0 (2 bits)
    reg [3:0] DirectionLights = 3'b000; // Directional lights (not fully utilized in this code)

    wire FlashFreq;  // Flash frequency generated by Adjust_Clk (slower clock signal)
    reg isFlash = 0;  // Flash control signal (1 bit) to enable or disable flashing

    // Instantiate Adjust_Clk to generate FlashFreq from the 50 MHz clock input
    Adjust_Clk c1(CLK_50MHz, FlashFreq);

    // Always block triggered on every rising edge of the 50 MHz clock (CLK_50MHz)
    always @(posedge CLK_50MHz) begin
        // Handle the idle state of the elevator when no floor is selected
        // The system enters calibration mode when it is at the initial state (floor 0)
        if (SelectedLevel == 2'b00 && CurrentLevel == 2'b00) begin
            UpPin <= 1'b0;    // Set UpPin to 0 (indicating the elevator is not moving up)
            DownPin <= 1'b1;  // Set DownPin to 1 (indicating the elevator is moving down)

            // Flashing LED pattern to indicate calibration mode
            if (FlashFreq) begin
                LevelLights <= 7'b00000000;  // Turn off all LEDs during one cycle of flashing
            end else begin
                LevelLights <= 7'b11111111;  // Turn on all LEDs during the next cycle of flashing
            end 

            // Floor switch handling: Update current and selected levels based on the active floor switch
            if (floorSwitch1) begin
                CurrentLevel <= 2'b01;  // Elevator is at floor 1
                SelectedLevel <= 2'b01;  // User has selected floor 1
                LevelLights <= 7'b1111001;  // LED pattern for floor 1
            end else if (floorSwitch2) begin
                CurrentLevel <= 2'b10;  // Elevator is at floor 2
                SelectedLevel <= 2'b10;  // User has selected floor 2
                LevelLights <= 7'b0100100;  // LED pattern for floor 2
            end else if (floorSwitch3) begin
                CurrentLevel <= 2'b11;  // Elevator is at floor 3
                SelectedLevel <= 2'b11;  // User has selected floor 3
                LevelLights <= 7'b0110000;  // LED pattern for floor 3
            end
            
            // Update each LED based on the current floor's LED pattern
            LEDA <= LevelLights[0];
            LEDB <= LevelLights[1];
            LEDC <= LevelLights[2];
            LEDD <= LevelLights[3];
            LEDE <= LevelLights[4];
            LEDF <= LevelLights[5];
            LEDG <= LevelLights[6];
        end else begin
            // When the elevator is not at the starting position, handle button presses for floor selection
            if (UpPin == 1'b0 && DownPin == 1'b0) begin
                // Check if any floor button is pressed (floorBtn1, floorBtn2, floorBtn3)
                if (floorBtn1) begin
                    SelectedLevel <= 2'b01;  // Select floor 1
                    LevelLights <= 7'b1111001;  // LED pattern for floor 1
                end
                else if (floorBtn2) begin
                    SelectedLevel <= 2'b10;  // Select floor 2
                    LevelLights <= 7'b0100100;  // LED pattern for floor 2
                end
                else if (floorBtn3) begin
                    SelectedLevel <= 2'b11;  // Select floor 3
                    LevelLights <= 7'b0110000;  // LED pattern for floor 3
                end
            end
            
            // Update the current floor based on the floor switch status (reed switches)
            if (floorSwitch1) begin
                CurrentLevel <= 2'b01;  // Elevator is at floor 1
            end else if (floorSwitch2) begin
                CurrentLevel <= 2'b10;  // Elevator is at floor 2
            end else if (floorSwitch3) begin
                CurrentLevel <= 2'b11;  // Elevator is at floor 3
            end 

            // Control the elevator movement direction based on selected and current levels
            if (SelectedLevel > CurrentLevel) begin
                UpPin <= 1'b1;    // Move elevator up
                DownPin <= 1'b0;  // Do not move down
            end else if (SelectedLevel < CurrentLevel) begin
                UpPin <= 1'b0;    // Do not move up
                DownPin <= 1'b1;  // Move elevator down
            end else begin
                UpPin <= 1'b0;    // Do not move (elevator is already at the correct floor)
                DownPin <= 1'b0;  // Do not move
            end
            
            // Set the flash condition if either up or down direction is active
            if ((UpPin == 1'b1 || DownPin == 1'b1)) begin
                isFlash = 1;  // Enable flashing when elevator is moving
            end else begin
                isFlash = 0;  // Disable flashing when elevator is idle
            end

            // If flashing is active and FlashFreq is true, blink the LEDs
            if (FlashFreq && isFlash) begin
                // Set all LEDs to high (off) for flashing effect
                LEDA <= 1'b1;
                LEDB <= 1'b1;
                LEDC <= 1'b1;
                LEDD <= 1'b1;
                LEDE <= 1'b1;
                LEDF <= 1'b1;
                LEDG <= 1'b1;
            end else begin
                // Otherwise, assign the current floor's LED pattern to each LED
                LEDA <= LevelLights[0];
                LEDB <= LevelLights[1];
                LEDC <= LevelLights[2];
                LEDD <= LevelLights[3];
                LEDE <= LevelLights[4];
                LEDF <= LevelLights[5];
                LEDG <= LevelLights[6];
            end
        end
    end
endmodule
